module ALU_tb;
	reg [31:0]A,B;
	reg [5:0] ALUFun;
	reg Sign;
	wire [31:0]S;
	
	ALU DUT(A,B,ALUFun,Sign,S);
	
	initial begin
		A=32'b1000_0000_0000_0000_0000_0000_0001_1111;
		B=32'b1111_1111_1111_1111_1111_0000_0000_0000;
		ALUFun=6'b000000;
		Sign=1;
 
		#200 ALUFun=6'b000001;
		#200 ALUFun=6'b011000;
		#200 ALUFun=6'b011110;
		#200 ALUFun=6'b010110;
		#200 ALUFun=6'b010001;
		#200 ALUFun=6'b011010;
		#200 ALUFun=6'b100000;
		#200 ALUFun=6'b100001;
		#200 ALUFun=6'b100011;
		#200 ALUFun=6'b110011;
		#200 ALUFun=6'b110001;
		#200 ALUFun=6'b110101;
		#200 ALUFun=6'b111101;
		#200 ALUFun=6'b111011;
		#200 ALUFun=6'b111111; 
		
		#200 Sign=0;
		
		#200 ALUFun=6'b000001;
		#200 ALUFun=6'b011000;
		#200 ALUFun=6'b011110;
		#200 ALUFun=6'b010110;
		#200 ALUFun=6'b010001;
		#200 ALUFun=6'b011010;
		#200 ALUFun=6'b100000;
		#200 ALUFun=6'b100001;
		#200 ALUFun=6'b100011;
		#200 ALUFun=6'b110011;
		#200 ALUFun=6'b110001;
		#200 ALUFun=6'b110101;
		#200 ALUFun=6'b111101;
		#200 ALUFun=6'b111011;
		#200 ALUFun=6'b111111; 
	end
endmodule